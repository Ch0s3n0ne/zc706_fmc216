-------------------------------------------------------------------------------------
-- FILE NAME : 
-- AUTHOR    : Luis
-- COMPANY   : 
-- UNITS     : Entity       - 
--             Architecture - Behavioral
-- LANGUAGE  : VHDL
-- DATE      : AUG 21, 2014
-------------------------------------------------------------------------------------
--
-------------------------------------------------------------------------------------
-- DESCRIPTION
-- ===========
-- 
-- 
-------------------------------------------------------------------------------------
 
-------------------------------------------------------------------------------------
-- LIBRARIES
-------------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_misc.all;
    use ieee.std_logic_arith.all; 

-------------------------------------------------------------------------------------
-- ENTITY
-------------------------------------------------------------------------------------
entity div_clock is
generic (
    TAP     : integer := 1
);
port (
    rst_in  : in  std_logic;
    clk_in  : in  std_logic;
    clk_out : out std_logic
);
end div_clock;

-------------------------------------------------------------------------------------
-- ARCHITECTURE
-------------------------------------------------------------------------------------
architecture Behavioral of div_clock is

-------------------------------------------------------------------------------------
-- CONSTANTS
-------------------------------------------------------------------------------------

-------------------------------------------------------------------------------------
-- SIGNALS
-------------------------------------------------------------------------------------
signal div_cnt : std_logic_vector(31 downto 0) := (others=>'0');

--***********************************************************************************
begin
--***********************************************************************************

process (clk_in, rst_in)
begin
   if rising_edge(clk_in) then
      if rst_in = '1' then
         div_cnt      <= (others=>'0');
         clk_out      <= '0';
      else 
         div_cnt <= div_cnt + 1;
         clk_out <= div_cnt(TAP);
      end if;
   end if;
end process;

--***********************************************************************************
end architecture Behavioral;
--***********************************************************************************

