-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : xcvr_fmc216_multi_gt.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module xcvr_fmc216_multi_gt (a Multi GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity xcvr_fmc216_multi_gt is
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "FALSE";        -- Set to "TRUE" to speed up sim reset
    RX_DFE_KL_CFG2_IN               : bit_vector :=  X"301148AC";
 
    PMA_RSV_IN                      : bit_vector :=  x"001E7080"
);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y20)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtnorthrefclk0_in                   : in   std_logic;
    gt0_gtnorthrefclk1_in                   : in   std_logic;
    gt0_gtsouthrefclk0_in                   : in   std_logic;
    gt0_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt0_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxdfelpmreset_in                    : in   std_logic;
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    gt0_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gtxtxn_out                          : out  std_logic;
    gt0_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;

    --GT1  (X0Y21)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtnorthrefclk0_in                   : in   std_logic;
    gt1_gtnorthrefclk1_in                   : in   std_logic;
    gt1_gtsouthrefclk0_in                   : in   std_logic;
    gt1_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt1_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxdfelpmreset_in                    : in   std_logic;
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    gt1_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gtxtxn_out                          : out  std_logic;
    gt1_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;

    --GT2  (X0Y22)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtnorthrefclk0_in                   : in   std_logic;
    gt2_gtnorthrefclk1_in                   : in   std_logic;
    gt2_gtsouthrefclk0_in                   : in   std_logic;
    gt2_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt2_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxdfelpmreset_in                    : in   std_logic;
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    gt2_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gtxtxn_out                          : out  std_logic;
    gt2_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;

    --GT3  (X0Y23)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtnorthrefclk0_in                   : in   std_logic;
    gt3_gtnorthrefclk1_in                   : in   std_logic;
    gt3_gtsouthrefclk0_in                   : in   std_logic;
    gt3_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt3_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxdfelpmreset_in                    : in   std_logic;
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    gt3_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gtxtxn_out                          : out  std_logic;
    gt3_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;

    --GT4  (X0Y24)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt4_gtnorthrefclk0_in                   : in   std_logic;
    gt4_gtnorthrefclk1_in                   : in   std_logic;
    gt4_gtsouthrefclk0_in                   : in   std_logic;
    gt4_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt4_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt4_rxlpmhfhold_in                      : in   std_logic;
    gt4_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxdfelpmreset_in                    : in   std_logic;
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    gt4_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    gt4_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt4_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt4_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gtxtxn_out                          : out  std_logic;
    gt4_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt4_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;

    --GT5  (X0Y25)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt5_gtnorthrefclk0_in                   : in   std_logic;
    gt5_gtnorthrefclk1_in                   : in   std_logic;
    gt5_gtsouthrefclk0_in                   : in   std_logic;
    gt5_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt5_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt5_rxlpmhfhold_in                      : in   std_logic;
    gt5_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxdfelpmreset_in                    : in   std_logic;
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    gt5_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    gt5_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt5_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt5_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gtxtxn_out                          : out  std_logic;
    gt5_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt5_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;

    --GT6  (X0Y26)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt6_gtnorthrefclk0_in                   : in   std_logic;
    gt6_gtnorthrefclk1_in                   : in   std_logic;
    gt6_gtsouthrefclk0_in                   : in   std_logic;
    gt6_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt6_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt6_rxlpmhfhold_in                      : in   std_logic;
    gt6_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxdfelpmreset_in                    : in   std_logic;
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    gt6_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    gt6_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt6_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt6_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gtxtxn_out                          : out  std_logic;
    gt6_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt6_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;

    --GT7  (X0Y27)
    --____________________________CHANNEL PORTS________________________________
    -------------------------- Channel - Clocking Ports ------------------------
    gt7_gtnorthrefclk0_in                   : in   std_logic;
    gt7_gtnorthrefclk1_in                   : in   std_logic;
    gt7_gtsouthrefclk0_in                   : in   std_logic;
    gt7_gtsouthrefclk1_in                   : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt7_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gtxrxn_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt7_rxlpmhfhold_in                      : in   std_logic;
    gt7_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxdfelpmreset_in                    : in   std_logic;
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    gt7_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    gt7_rxpmareset_in                       : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    gt7_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt7_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gtxtxn_out                          : out  std_logic;
    gt7_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt7_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;


    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN : in std_logic;
     GT0_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT1_QPLLOUTCLK_IN : in std_logic;
     GT1_QPLLOUTREFCLK_IN : in std_logic

);


end xcvr_fmc216_multi_gt;
    
architecture RTL of xcvr_fmc216_multi_gt is
    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "xcvr_fmc216_multi_gt,gtwizard_v3_6_13,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;
    signal   gt0_qplloutclk_i         :   std_logic;
    signal   gt0_qplloutrefclk_i      :   std_logic;
    signal   gt1_qplloutclk_i         :   std_logic;
    signal   gt1_qplloutrefclk_i      :   std_logic;

    signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt4_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt4_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt5_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt5_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt6_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt6_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
    signal  gt7_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt7_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
    signal   gt0_qpllclk_i            :   std_logic;
    signal   gt0_qpllrefclk_i         :   std_logic;
    signal   gt1_qpllclk_i            :   std_logic;
    signal   gt1_qpllrefclk_i         :   std_logic;
    signal   gt2_qpllclk_i            :   std_logic;
    signal   gt2_qpllrefclk_i         :   std_logic;
    signal   gt3_qpllclk_i            :   std_logic;
    signal   gt3_qpllrefclk_i         :   std_logic;
    signal   gt4_qpllclk_i            :   std_logic;
    signal   gt4_qpllrefclk_i         :   std_logic;
    signal   gt5_qpllclk_i            :   std_logic;
    signal   gt5_qpllrefclk_i         :   std_logic;
    signal   gt6_qpllclk_i            :   std_logic;
    signal   gt6_qpllrefclk_i         :   std_logic;
    signal   gt7_qpllclk_i            :   std_logic;
    signal   gt7_qpllrefclk_i         :   std_logic;
    signal   gt0_cpllreset_i            :   std_logic;
    signal   gt0_cpllpd_i         :   std_logic;
    signal   gt1_cpllreset_i            :   std_logic;
    signal   gt1_cpllpd_i         :   std_logic;
    signal   gt2_cpllreset_i            :   std_logic;
    signal   gt2_cpllpd_i         :   std_logic;
    signal   gt3_cpllreset_i            :   std_logic;
    signal   gt3_cpllpd_i         :   std_logic;
    signal   gt4_cpllreset_i            :   std_logic;
    signal   gt4_cpllpd_i         :   std_logic;
    signal   gt5_cpllreset_i            :   std_logic;
    signal   gt5_cpllpd_i         :   std_logic;
    signal   gt6_cpllreset_i            :   std_logic;
    signal   gt6_cpllpd_i         :   std_logic;
    signal   gt7_cpllreset_i            :   std_logic;
    signal   gt7_cpllpd_i         :   std_logic;

--*************************** Component Declarations **************************
component xcvr_fmc216_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP       : string   := "FALSE";
    RX_DFE_KL_CFG2_IN            : bit_vector :=   X"3010D90C";
    PMA_RSV_IN                   : bit_vector :=   X"00000000";
    SIM_CPLLREFCLK_SEL           : bit_vector :=   "001";
    PCS_RSVD_ATTR_IN             : bit_vector :=   X"000000000000"
);
port 
(   
     cpllrefclksel_in : in std_logic_vector (2 downto 0);
    -------------------------- Channel - Clocking Ports ------------------------
    gtnorthrefclk0_in                       : in   std_logic;
    gtnorthrefclk1_in                       : in   std_logic;
    gtsouthrefclk0_in                       : in   std_logic;
    gtsouthrefclk1_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    drpaddr_in                              : in   std_logic_vector(8 downto 0);
    drpclk_in                               : in   std_logic;
    drpdi_in                                : in   std_logic_vector(15 downto 0);
    drpdo_out                               : out  std_logic_vector(15 downto 0);
    drpen_in                                : in   std_logic;
    drprdy_out                              : out  std_logic;
    drpwe_in                                : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    qpllclk_in                              : in   std_logic;
    qpllrefclk_in                           : in   std_logic;
    --------------------------- Digital Monitor Ports --------------------------
    dmonitorout_out                         : out  std_logic_vector(7 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    eyescanreset_in                         : in   std_logic;
    rxuserrdy_in                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    eyescandataerror_out                    : out  std_logic;
    eyescantrigger_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    rxusrclk_in                             : in   std_logic;
    rxusrclk2_in                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    rxdata_out                              : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    rxdisperr_out                           : out  std_logic_vector(3 downto 0);
    rxnotintable_out                        : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gtxrxp_in                               : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gtxrxn_in                               : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    rxlpmhfhold_in                          : in   std_logic;
    rxlpmlfhold_in                          : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    rxdfelpmreset_in                        : in   std_logic;
    rxmonitorout_out                        : out  std_logic_vector(6 downto 0);
    rxmonitorsel_in                         : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    rxoutclk_out                            : out  std_logic;
    rxoutclkfabric_out                      : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gtrxreset_in                            : in   std_logic;
    rxpmareset_in                           : in   std_logic;
    ---------------------- Receive Ports - RX gearbox ports --------------------
    rxslide_in                              : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    rxchariscomma_out                       : out  std_logic_vector(3 downto 0);
    rxcharisk_out                           : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    rxresetdone_out                         : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gttxreset_in                            : in   std_logic;
    txuserrdy_in                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    txusrclk_in                             : in   std_logic;
    txusrclk2_in                            : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    txdata_in                               : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gtxtxn_out                              : out  std_logic;
    gtxtxp_out                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    txoutclk_out                            : out  std_logic;
    txoutclkfabric_out                      : out  std_logic;
    txoutclkpcs_out                         : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    txcharisk_in                            : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    txresetdone_out                         : out  std_logic


);
end component;



--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt0_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 

    gt1_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt1_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 

    gt2_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt2_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 

    gt3_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt3_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 

    gt4_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt4_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 

    gt5_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt5_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 

    gt6_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt6_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 

    gt7_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt7_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 


 
    --------------------------- GT Instances  -------------------------------   
 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y20)

gt0_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt0_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt0_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt0_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt0_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt0_drpaddr_in,
        drpclk_in                       =>      gt0_drpclk_in,
        drpdi_in                        =>      gt0_drpdi_in,
        drpdo_out                       =>      gt0_drpdo_out,
        drpen_in                        =>      gt0_drpen_in,
        drprdy_out                      =>      gt0_drprdy_out,
        drpwe_in                        =>      gt0_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt0_qpllclk_i,
        qpllrefclk_in                   =>      gt0_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt0_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt0_eyescanreset_in,
        rxuserrdy_in                    =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt0_eyescandataerror_out,
        eyescantrigger_in               =>      gt0_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt0_rxusrclk_in,
        rxusrclk2_in                    =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt0_rxdisperr_out,
        rxnotintable_out                =>      gt0_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt0_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt0_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt0_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt0_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt0_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt0_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt0_rxoutclk_out,
        rxoutclkfabric_out              =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt0_gtrxreset_in,
        rxpmareset_in                   =>      gt0_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt0_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt0_rxchariscomma_out,
        rxcharisk_out                   =>      gt0_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt0_gttxreset_in,
        txuserrdy_in                    =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt0_txusrclk_in,
        txusrclk2_in                    =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt0_gtxtxn_out,
        gtxtxp_out                      =>      gt0_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt0_txoutclk_out,
        txoutclkfabric_out              =>      gt0_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt0_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt0_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt0_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y21)

gt1_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt1_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt1_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt1_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt1_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt1_drpaddr_in,
        drpclk_in                       =>      gt1_drpclk_in,
        drpdi_in                        =>      gt1_drpdi_in,
        drpdo_out                       =>      gt1_drpdo_out,
        drpen_in                        =>      gt1_drpen_in,
        drprdy_out                      =>      gt1_drprdy_out,
        drpwe_in                        =>      gt1_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt1_qpllclk_i,
        qpllrefclk_in                   =>      gt1_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt1_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt1_eyescanreset_in,
        rxuserrdy_in                    =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt1_eyescandataerror_out,
        eyescantrigger_in               =>      gt1_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt1_rxusrclk_in,
        rxusrclk2_in                    =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt1_rxdisperr_out,
        rxnotintable_out                =>      gt1_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt1_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt1_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt1_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt1_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt1_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt1_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt1_rxoutclk_out,
        rxoutclkfabric_out              =>      gt1_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt1_gtrxreset_in,
        rxpmareset_in                   =>      gt1_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt1_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt1_rxchariscomma_out,
        rxcharisk_out                   =>      gt1_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt1_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt1_gttxreset_in,
        txuserrdy_in                    =>      gt1_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt1_txusrclk_in,
        txusrclk2_in                    =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt1_gtxtxn_out,
        gtxtxp_out                      =>      gt1_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt1_txoutclk_out,
        txoutclkfabric_out              =>      gt1_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt1_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt1_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt1_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y22)

gt2_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt2_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt2_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt2_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt2_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt2_drpaddr_in,
        drpclk_in                       =>      gt2_drpclk_in,
        drpdi_in                        =>      gt2_drpdi_in,
        drpdo_out                       =>      gt2_drpdo_out,
        drpen_in                        =>      gt2_drpen_in,
        drprdy_out                      =>      gt2_drprdy_out,
        drpwe_in                        =>      gt2_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt2_qpllclk_i,
        qpllrefclk_in                   =>      gt2_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt2_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt2_eyescanreset_in,
        rxuserrdy_in                    =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt2_eyescandataerror_out,
        eyescantrigger_in               =>      gt2_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt2_rxusrclk_in,
        rxusrclk2_in                    =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt2_rxdisperr_out,
        rxnotintable_out                =>      gt2_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt2_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt2_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt2_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt2_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt2_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt2_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt2_rxoutclk_out,
        rxoutclkfabric_out              =>      gt2_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt2_gtrxreset_in,
        rxpmareset_in                   =>      gt2_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt2_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt2_rxchariscomma_out,
        rxcharisk_out                   =>      gt2_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt2_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt2_gttxreset_in,
        txuserrdy_in                    =>      gt2_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt2_txusrclk_in,
        txusrclk2_in                    =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt2_gtxtxn_out,
        gtxtxp_out                      =>      gt2_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt2_txoutclk_out,
        txoutclkfabric_out              =>      gt2_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt2_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt2_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt2_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y23)

gt3_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt3_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt3_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt3_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt3_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt3_drpaddr_in,
        drpclk_in                       =>      gt3_drpclk_in,
        drpdi_in                        =>      gt3_drpdi_in,
        drpdo_out                       =>      gt3_drpdo_out,
        drpen_in                        =>      gt3_drpen_in,
        drprdy_out                      =>      gt3_drprdy_out,
        drpwe_in                        =>      gt3_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt3_qpllclk_i,
        qpllrefclk_in                   =>      gt3_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt3_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt3_eyescanreset_in,
        rxuserrdy_in                    =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt3_eyescandataerror_out,
        eyescantrigger_in               =>      gt3_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt3_rxusrclk_in,
        rxusrclk2_in                    =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt3_rxdisperr_out,
        rxnotintable_out                =>      gt3_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt3_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt3_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt3_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt3_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt3_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt3_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt3_rxoutclk_out,
        rxoutclkfabric_out              =>      gt3_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt3_gtrxreset_in,
        rxpmareset_in                   =>      gt3_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt3_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt3_rxchariscomma_out,
        rxcharisk_out                   =>      gt3_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt3_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt3_gttxreset_in,
        txuserrdy_in                    =>      gt3_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt3_txusrclk_in,
        txusrclk2_in                    =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt3_gtxtxn_out,
        gtxtxp_out                      =>      gt3_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt3_txoutclk_out,
        txoutclkfabric_out              =>      gt3_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt3_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt3_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt3_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT4  (X0Y24)

gt4_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt4_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt4_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt4_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt4_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt4_drpaddr_in,
        drpclk_in                       =>      gt4_drpclk_in,
        drpdi_in                        =>      gt4_drpdi_in,
        drpdo_out                       =>      gt4_drpdo_out,
        drpen_in                        =>      gt4_drpen_in,
        drprdy_out                      =>      gt4_drprdy_out,
        drpwe_in                        =>      gt4_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt4_qpllclk_i,
        qpllrefclk_in                   =>      gt4_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt4_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt4_eyescanreset_in,
        rxuserrdy_in                    =>      gt4_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt4_eyescandataerror_out,
        eyescantrigger_in               =>      gt4_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt4_rxusrclk_in,
        rxusrclk2_in                    =>      gt4_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt4_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt4_rxdisperr_out,
        rxnotintable_out                =>      gt4_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt4_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt4_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt4_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt4_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt4_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt4_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt4_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt4_rxoutclk_out,
        rxoutclkfabric_out              =>      gt4_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt4_gtrxreset_in,
        rxpmareset_in                   =>      gt4_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt4_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt4_rxchariscomma_out,
        rxcharisk_out                   =>      gt4_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt4_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt4_gttxreset_in,
        txuserrdy_in                    =>      gt4_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt4_txusrclk_in,
        txusrclk2_in                    =>      gt4_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt4_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt4_gtxtxn_out,
        gtxtxp_out                      =>      gt4_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt4_txoutclk_out,
        txoutclkfabric_out              =>      gt4_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt4_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt4_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt4_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT5  (X0Y25)

gt5_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt5_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt5_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt5_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt5_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt5_drpaddr_in,
        drpclk_in                       =>      gt5_drpclk_in,
        drpdi_in                        =>      gt5_drpdi_in,
        drpdo_out                       =>      gt5_drpdo_out,
        drpen_in                        =>      gt5_drpen_in,
        drprdy_out                      =>      gt5_drprdy_out,
        drpwe_in                        =>      gt5_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt5_qpllclk_i,
        qpllrefclk_in                   =>      gt5_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt5_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt5_eyescanreset_in,
        rxuserrdy_in                    =>      gt5_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt5_eyescandataerror_out,
        eyescantrigger_in               =>      gt5_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt5_rxusrclk_in,
        rxusrclk2_in                    =>      gt5_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt5_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt5_rxdisperr_out,
        rxnotintable_out                =>      gt5_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt5_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt5_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt5_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt5_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt5_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt5_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt5_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt5_rxoutclk_out,
        rxoutclkfabric_out              =>      gt5_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt5_gtrxreset_in,
        rxpmareset_in                   =>      gt5_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt5_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt5_rxchariscomma_out,
        rxcharisk_out                   =>      gt5_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt5_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt5_gttxreset_in,
        txuserrdy_in                    =>      gt5_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt5_txusrclk_in,
        txusrclk2_in                    =>      gt5_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt5_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt5_gtxtxn_out,
        gtxtxp_out                      =>      gt5_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt5_txoutclk_out,
        txoutclkfabric_out              =>      gt5_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt5_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt5_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt5_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT6  (X0Y26)

gt6_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt6_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt6_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt6_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt6_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt6_drpaddr_in,
        drpclk_in                       =>      gt6_drpclk_in,
        drpdi_in                        =>      gt6_drpdi_in,
        drpdo_out                       =>      gt6_drpdo_out,
        drpen_in                        =>      gt6_drpen_in,
        drprdy_out                      =>      gt6_drprdy_out,
        drpwe_in                        =>      gt6_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt6_qpllclk_i,
        qpllrefclk_in                   =>      gt6_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt6_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt6_eyescanreset_in,
        rxuserrdy_in                    =>      gt6_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt6_eyescandataerror_out,
        eyescantrigger_in               =>      gt6_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt6_rxusrclk_in,
        rxusrclk2_in                    =>      gt6_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt6_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt6_rxdisperr_out,
        rxnotintable_out                =>      gt6_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt6_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt6_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt6_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt6_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt6_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt6_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt6_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt6_rxoutclk_out,
        rxoutclkfabric_out              =>      gt6_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt6_gtrxreset_in,
        rxpmareset_in                   =>      gt6_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt6_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt6_rxchariscomma_out,
        rxcharisk_out                   =>      gt6_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt6_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt6_gttxreset_in,
        txuserrdy_in                    =>      gt6_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt6_txusrclk_in,
        txusrclk2_in                    =>      gt6_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt6_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt6_gtxtxn_out,
        gtxtxp_out                      =>      gt6_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt6_txoutclk_out,
        txoutclkfabric_out              =>      gt6_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt6_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt6_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt6_txresetdone_out

    );

 

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT7  (X0Y27)

gt7_xcvr_fmc216_i : xcvr_fmc216_GT 
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        SIM_CPLLREFCLK_SEL            =>  "001",
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        cpllrefclksel_in => "001",
        -------------------------- Channel - Clocking Ports ------------------------
        gtnorthrefclk0_in               =>      gt7_gtnorthrefclk0_in,
        gtnorthrefclk1_in               =>      gt7_gtnorthrefclk1_in,
        gtsouthrefclk0_in               =>      gt7_gtsouthrefclk0_in,
        gtsouthrefclk1_in               =>      gt7_gtsouthrefclk1_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt7_drpaddr_in,
        drpclk_in                       =>      gt7_drpclk_in,
        drpdi_in                        =>      gt7_drpdi_in,
        drpdo_out                       =>      gt7_drpdo_out,
        drpen_in                        =>      gt7_drpen_in,
        drprdy_out                      =>      gt7_drprdy_out,
        drpwe_in                        =>      gt7_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt7_qpllclk_i,
        qpllrefclk_in                   =>      gt7_qpllrefclk_i,
        --------------------------- Digital Monitor Ports --------------------------
        dmonitorout_out                 =>      gt7_dmonitorout_out,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt7_eyescanreset_in,
        rxuserrdy_in                    =>      gt7_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt7_eyescandataerror_out,
        eyescantrigger_in               =>      gt7_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt7_rxusrclk_in,
        rxusrclk2_in                    =>      gt7_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt7_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt7_rxdisperr_out,
        rxnotintable_out                =>      gt7_rxnotintable_out,
        --------------------------- Receive Ports - RX AFE -------------------------
        gtxrxp_in                       =>      gt7_gtxrxp_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtxrxn_in                       =>      gt7_gtxrxn_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt7_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt7_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfelpmreset_in                =>      gt7_rxdfelpmreset_in,
        rxmonitorout_out                =>      gt7_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt7_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt7_rxoutclk_out,
        rxoutclkfabric_out              =>      gt7_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt7_gtrxreset_in,
        rxpmareset_in                   =>      gt7_rxpmareset_in,
        ---------------------- Receive Ports - RX gearbox ports --------------------
        rxslide_in                      =>      gt7_rxslide_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxchariscomma_out               =>      gt7_rxchariscomma_out,
        rxcharisk_out                   =>      gt7_rxcharisk_out,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt7_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt7_gttxreset_in,
        txuserrdy_in                    =>      gt7_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt7_txusrclk_in,
        txusrclk2_in                    =>      gt7_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt7_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gtxtxn_out                      =>      gt7_gtxtxn_out,
        gtxtxp_out                      =>      gt7_gtxtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt7_txoutclk_out,
        txoutclkfabric_out              =>      gt7_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt7_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        txcharisk_in                    =>      gt7_txcharisk_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt7_txresetdone_out

    );


end RTL;     
